module data_memory(
    input logic clk, rst,
    input logic [31:0] A,
    input logic [31:0] WD,
    input logic WE,
    output logic [31:0] RD,
    output logic [31:0] prode
);
    
endmodule